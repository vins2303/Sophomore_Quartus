library verilog;
use verilog.vl_types.all;
entity Sort2_vlg_vec_tst is
end Sort2_vlg_vec_tst;
