library verilog;
use verilog.vl_types.all;
entity N2_vlg_vec_tst is
end N2_vlg_vec_tst;
