library verilog;
use verilog.vl_types.all;
entity N4_vlg_vec_tst is
end N4_vlg_vec_tst;
