library verilog;
use verilog.vl_types.all;
entity Sort2_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        in_data         : in     vl_logic_vector(7 downto 0);
        isData          : in     vl_logic;
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Sort2_vlg_sample_tst;
