library verilog;
use verilog.vl_types.all;
entity N1_vlg_vec_tst is
end N1_vlg_vec_tst;
