library verilog;
use verilog.vl_types.all;
entity sort3_vlg_vec_tst is
end sort3_vlg_vec_tst;
