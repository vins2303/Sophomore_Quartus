library verilog;
use verilog.vl_types.all;
entity cyclonev_and1 is
    port(
        Y               : out    vl_logic;
        IN1             : in     vl_logic
    );
end cyclonev_and1;
