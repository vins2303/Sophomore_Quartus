library verilog;
use verilog.vl_types.all;
entity N3_vlg_vec_tst is
end N3_vlg_vec_tst;
