library verilog;
use verilog.vl_types.all;
entity N2 is
    port(
        clk             : in     vl_logic;
        \in\            : in     vl_logic;
        \out\           : out    vl_logic;
        rst             : in     vl_logic
    );
end N2;
