`include "Module/Roles.v"
`include "Module/Cactus.v"
`include "Module/VGA.v"
`include "Module/IR_RECEIVE.V"
`include "Module/BCD_16bit.v"
`include "Module/Segment_7.v"
module End(
	input clk, rst,		//clk 50MHz
	input Stop_SW,
	output  VGA_HS, VGA_VS,
	output reg [7:0] VGA_R,VGA_G,VGA_B,
	output VGA_BLANK_N,VGA_CLOCK,
	input IRDA_RXD,
	output [4:0] Speed_Led,
	output [6:0] HEX0, HEX1, HEX2, HEX3
);
	wire Game_rst = rst && (IR_Pos_Ready == 1 && IR_Ready == 0 && IR_data[23:16] == 8'h12) ? 0 : 1;

	/*----------------------------- Clk ---------------------------------------*/
	reg clk25M;
	always@(posedge clk) clk25M = ~clk25M;
	reg clk_1K; // 0.001s
	reg clk_500;
	reg clk_250;
	reg clk_125;
	reg clk_62;
	reg clk_31;
	reg clk_15;
	reg clk_7;
	reg clk_3;
	reg clk_1;
	reg [21:0]clk_1K_count;
	
	always@(posedge clk_1K ) clk_500 <= ~clk_500;
	always@(posedge clk_500) clk_250 <= ~clk_250;
	always@(posedge clk_250) clk_125 <= ~clk_125;
	always@(posedge clk_125) clk_62  <= ~clk_62;
	always@(posedge clk_62 ) clk_31  <= ~clk_31;
	always@(posedge clk_31 ) clk_15  <= ~clk_15;
	always@(posedge clk_15 ) clk_7   <= ~clk_7;
	always@(posedge clk_7  ) clk_3   <= ~clk_3;
	always@(posedge clk_3  ) clk_1   <= ~clk_1;

	always@(posedge clk, negedge rst)begin
		if(!rst) begin
			clk_1K_count <= 0;
		end else begin
			if(clk_1K_count < 25000)
				clk_1K_count <= clk_1K_count + 1;
			else begin
				clk_1K_count <= 0;
				clk_1K <= ~clk_1K;
			end 

		end
	end
	/*----------------------------------- VGA --------------------------------------*/
	wire [12:0] VGA_X,VGA_Y;

	VGA vga_
	(
		.clk25M(clk25M),
		.rst(rst),
		.VGA_HS(VGA_HS),
		.VGA_VS(VGA_VS),
		.VGA_BLANK_N(VGA_BLANK_N), 
		.VGA_CLOCK(VGA_CLOCK), 
		.X(VGA_X), 
		.Y(VGA_Y)
	);

	always@(posedge clk25M) begin
		if (!rst) begin
			{VGA_R,VGA_G,VGA_B}<=0;
		end else 
		begin
			if(Game_Stop) begin
				if(VGA_X < 276 && VGA_Y < 86)
					{VGA_R,VGA_G,VGA_B} <= Ranther_Image[VGA_Y][ VGA_X] ? 24'h00FFFF : Back_Color;
				else
					{VGA_R,VGA_G,VGA_B} <= Back_Color;

			end else begin
				if((VGA_X < Roles_Point_X + Roles_Width && VGA_X >= Roles_Point_X) && (VGA_Y < Roles_Point_Y + Roles_Heigh && VGA_Y >= Roles_Point_Y)) begin
					{VGA_R,VGA_G,VGA_B} <= ( Roles_Image_Status ? Roles_Image_1[VGA_Y - Roles_Point_Y][ VGA_X - Roles_Point_X] : Roles_Image_2[VGA_Y - Roles_Point_Y][ VGA_X - Roles_Point_X] ) ? Roles_Color :24'h000000;

				end else if((VGA_X < Roles_Fire_Point_X + Roles_Fire_Width && VGA_X >= Roles_Fire_Point_X) && (VGA_Y < Roles_Fire_Point_Y + Roles_Fire_Heigh && VGA_Y >= Roles_Fire_Point_Y)) begin
					{VGA_R,VGA_G,VGA_B} <= Fire_Image[VGA_Y - Roles_Fire_Point_Y][ VGA_X - Roles_Fire_Point_X] ? Fire_Color : Back_Color;

				end else if((VGA_X < Cactus_Point_X_0 + Cactus_Width_0 && VGA_X >= Cactus_Point_X_0) && (VGA_Y < Cactus_Point_Y_0 + Cactus_Heigh_0 && VGA_Y >= Cactus_Point_Y_0)) begin
					{VGA_R,VGA_G,VGA_B} <= Cactus_Image[VGA_Y - Cactus_Point_Y_0][ VGA_X - Cactus_Point_X_0] ? Cactus_Color : Back_Color;

				end else if(VGA_Y == 400) begin
					{VGA_R,VGA_G,VGA_B} <= Floor_Color;

				end else begin
					{VGA_R,VGA_G,VGA_B} <= Back_Color;

				end
			end
		end
	end
/*------------------------------- Color ---------------------------------*/
	parameter Roles_Color  = 24'h91f0fa;
	parameter Cactus_Color = 24'h94fda2;
	parameter Back_Color   = 24'h000000;
	parameter Floor_Color  = 24'h048787;
	parameter Fire_Color   = 24'hFF3333;

/*------------------------------ IR ----------------------------------------*/
	wire [31:0] IR_data;
	wire IR_Ready;
	reg  IR_Pos_Ready;
	IR_RECEIVE IR_1(clk,rst,IRDA_RXD,IR_Ready,IR_data);
	always@(posedge clk) IR_Pos_Ready <= IR_Ready;

/*------------------------------ Game_Start --------------------------------*/
	reg Game_Start;
	always@(negedge Game_rst, negedge IR_Ready) begin
		if(!Game_rst) 
			Game_Start <= 1;
		else if(IR_data[23:16] == 8'h16)
			Game_Start <= ~Game_Start;
	end

/* ----------------------------- Fraction ----------------------------- */
	reg [15:0] Game_Fraction;
	wire [15:0] Game_Fraction_BCD;
	BCD_16bit bcd_16bit(.bin( Game_Fraction), .out( Game_Fraction_BCD));
	Segment_7 hex_0(.num( Game_Fraction_BCD[3 : 0]), .out(HEX0));
	Segment_7 hex_1(.num( Game_Fraction_BCD[7 : 4]), .out(HEX1));
	Segment_7 hex_2(.num( Game_Fraction_BCD[11: 8]), .out(HEX2));
	Segment_7 hex_3(.num( Game_Fraction_BCD[15:12]), .out(HEX3));

	always@(posedge Cactus_clk, negedge Game_rst) begin
		if(!Game_rst) begin 
			Game_Fraction <= 0;
		end else begin
			if(Cactus_Point_X_0 < 1 && !Game_Stop) Game_Fraction <= Game_Fraction + 1;
		end
	end

/*------------------------------ Stop ---------------------------------------*/
	wire Game_Stop;
	assign Game_Stop = isOverlap_Stop || Stop_SW || Game_Start;

/*------------------------------ isOverlap--------------------------------*/
	reg isOverlap_Stop;
	always@(posedge clk, negedge Game_rst)begin
		if(!Game_rst)begin
			isOverlap_Stop <= 0;
			
		end else begin
			if((Roles_Point_X    + Roles_Width    > Cactus_Point_X_0   &&  
			    Cactus_Point_X_0 + Cactus_Width_0 > Roles_Point_X    ) &&
			   (Roles_Point_Y    + Roles_Heigh    > Cactus_Point_Y_0   && 
				Cactus_Point_Y_0 + Cactus_Heigh_0 > Roles_Point_Y  ))
			begin
				
				isOverlap_Stop <= 1;	
			end
		end
	end

/*----------------------------- Roles ----------------------------------*/
	wire Roles_Jump;

	parameter Roles_Width = 40;
	parameter Roles_Heigh = 43;

	wire [9:0] Roles_Point_X;
	wire [9:0] Roles_Point_Y;
	Roles #(Roles_Width, Roles_Heigh)  roles_
	(
		.clk(clk_31), 
		.rst(Game_rst), 
		.Stop(Game_Stop),
		.Point_X( Roles_Point_X), 
		.Point_Y( Roles_Point_Y),
		.Jump_Button(Roles_Jump)
	);

/*----------------------------- Roles_Jump ----------------------------------*/
	assign Roles_Jump = (IR_Pos_Ready == 1 && IR_Ready == 0 && IR_data[23:16] == 8'h1A) ? 1 : 0;

/*----------------------------- Roles_Fire ----------------------------------*/
	parameter Roles_Fire_Width = 18;
	parameter Roles_Fire_Heigh = 10;
	wire [9:0] Roles_Fire_Point_X;
	wire [9:0] Roles_Fire_Point_Y;

	assign Roles_Fire_Point_X = Roles_Point_X + Roles_Width + 5;
	assign Roles_Fire_Point_Y = Roles_Fire_Run ? Roles_Point_Y + 13 : 1000;

	reg Roles_Fire_Run;
	reg pos_clk_1;

	always@(posedge clk) pos_clk_1 <= clk_1;

	always@(posedge clk, negedge Game_rst) begin
		if(!Game_rst) begin
			Roles_Fire_Run <= 0;
		end else begin
			if(IR_Pos_Ready == 1 && IR_Ready == 0 && IR_data[23:16] == 8'h01 && !Game_Stop) begin
				Roles_Fire_Run <= 1;
			end else if(Roles_Fire_Run == 1 && pos_clk_1 == 0 && clk_1 == 1) begin
				Roles_Fire_Run <= 0;
			end
		end
	end

/*----------------------------- Cactus Speed ---------------------------------*/
	reg Cactus_clk;
	reg [3:0] Game_Speed;
	always@(negedge IR_Ready,negedge Game_rst)begin
		if(Game_rst == 0)begin
			Game_Speed <= 2;
		end else begin
			case(IR_data[23:16])
				8'h1B: if(Game_Speed < 5) Game_Speed <= Game_Speed + 1;
				8'h1F: if(Game_Speed > 0) Game_Speed <= Game_Speed - 1;

				default:;
			endcase
		end
	end


	always@(posedge clk) begin
		case(Game_Speed)
			0: Cactus_clk <= clk_31;
			1: Cactus_clk <= clk_62;
			2: Cactus_clk <= clk_125;
			3: Cactus_clk <= clk_250;
			4: Cactus_clk <= clk_250;
			5: Cactus_clk <= clk_500;
			default: Cactus_clk <= clk;
		endcase
	end

	assign Speed_Led[0] = Game_Speed>0;
	assign Speed_Led[1] = Game_Speed>1;
	assign Speed_Led[2] = Game_Speed>2;
	assign Speed_Led[3] = Game_Speed>3;
	assign Speed_Led[4] = Game_Speed>4;

/*----------------------------- Cactus ---------------------------------*/
	wire [9:0] Cactus_Point_X_0;
	wire [9:0] Cactus_Point_Y_0;
	parameter Cactus_Width_0 = 15;
	parameter Cactus_Heigh_0 = 33;
	reg Cactus_Wipe_0;

	Cactus #(Cactus_Width_0, Cactus_Heigh_0) Cactus_ 
	(
		.clk(     Cactus_clk       ), 
		.rst(     Game_rst         ), 
		.Stop(    Game_Stop        ),
		.Point_X( Cactus_Point_X_0 ), 
		.Point_Y( Cactus_Point_Y_0 ),
		.Wipe(    Cactus_Wipe_0    )
	);


	always@(posedge clk, negedge Game_rst) begin
		if(!Game_rst) begin
			Cactus_Wipe_0 <= 0;
		end else begin
			if( (Roles_Fire_Point_X + Roles_Fire_Width > Cactus_Point_X_0     &&  
			     Cactus_Point_X_0   + Cactus_Width_0   > Roles_Fire_Point_X ) &&
				(Roles_Fire_Point_Y + Roles_Fire_Heigh > Cactus_Point_Y_0     && 
				 Cactus_Point_Y_0   + Cactus_Heigh_0   > Roles_Fire_Point_Y ) )
			begin
				Cactus_Wipe_0 <= 1;
			end else if(pos_clk_1 == 0 && clk_1 == 1 && Cactus_Wipe_0 == 1) begin 
				Cactus_Wipe_0 <= 0;
			end
		end
	end

/*------------------------------- Image -------------------------------*/
reg Roles_Image_Status;

always@(posedge clk_7) if(!Game_Stop) Roles_Image_Status <= ~Roles_Image_Status;

wire [ 0 : 39] Roles_Image_1[ 0 : 42];

assign Roles_Image_1[0] = 40'b0000000000000000000000111111111111111100;
assign Roles_Image_1[1] = 40'b0000000000000000000000111111111111111100;
assign Roles_Image_1[2] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[3] = 40'b0000000000000000000011110011111111111111;
assign Roles_Image_1[4] = 40'b0000000000000000000011110011111111111111;
assign Roles_Image_1[5] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[6] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[7] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[8] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[9] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[10] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_1[11] = 40'b0000000000000000000011111111110000000000;
assign Roles_Image_1[12] = 40'b0000000000000000000011111111110000000000;
assign Roles_Image_1[13] = 40'b0000000000000000000011111111111111110000;
assign Roles_Image_1[14] = 40'b0000000000000000000011111111111111110000;
assign Roles_Image_1[15] = 40'b1100000000000000001111111111000000000000;
assign Roles_Image_1[16] = 40'b1100000000000000001111111111000000000000;
assign Roles_Image_1[17] = 40'b1100000000000001111111111111000000000000;
assign Roles_Image_1[18] = 40'b1100000000000001111111111111000000000000;
assign Roles_Image_1[19] = 40'b1111000000001111111111111111111100000000;
assign Roles_Image_1[20] = 40'b1111000000001111111111111111111100000000;
assign Roles_Image_1[21] = 40'b1111110000111111111111111111001100000000;
assign Roles_Image_1[22] = 40'b1111110000111111111111111111001100000000;
assign Roles_Image_1[23] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_1[24] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_1[25] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_1[26] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_1[27] = 40'b0011111111111111111111111111000000000000;
assign Roles_Image_1[28] = 40'b0011111111111111111111111100000000000000;
assign Roles_Image_1[29] = 40'b0000111111111111111111111100000000000000;
assign Roles_Image_1[30] = 40'b0000111111111111111111111100000000000000;
assign Roles_Image_1[31] = 40'b0000001111111111111111110000000000000000;
assign Roles_Image_1[32] = 40'b0000001111111111111111110000000000000000;
assign Roles_Image_1[33] = 40'b0000000011111111111111000000000000000000;
assign Roles_Image_1[34] = 40'b0000000011111111111111000000000000000000;
assign Roles_Image_1[35] = 40'b0000000000111100001111000000000000000000;
assign Roles_Image_1[36] = 40'b0000000000111100001111000000000000000000;
assign Roles_Image_1[37] = 40'b0000000000001111000011000000000000000000;
assign Roles_Image_1[38] = 40'b0000000000001111000011000000000000000000;
assign Roles_Image_1[39] = 40'b0000000000000000000011000000000000000000;
assign Roles_Image_1[40] = 40'b0000000000000000000011000000000000000000;
assign Roles_Image_1[41] = 40'b0000000000000000000011110000000000000000;
assign Roles_Image_1[42] = 40'b0000000000000000000011110000000000000000;

wire [ 0 : 39] Roles_Image_2[ 0 : 42];
assign Roles_Image_2[0] = 40'b0000000000000000000000111111111111111100;
assign Roles_Image_2[1] = 40'b0000000000000000000000111111111111111100;
assign Roles_Image_2[2] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[3] = 40'b0000000000000000000011110011111111111111;
assign Roles_Image_2[4] = 40'b0000000000000000000011110011111111111111;
assign Roles_Image_2[5] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[6] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[7] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[8] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[9] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[10] = 40'b0000000000000000000011111111111111111111;
assign Roles_Image_2[11] = 40'b0000000000000000000011111111110000000000;
assign Roles_Image_2[12] = 40'b0000000000000000000011111111110000000000;
assign Roles_Image_2[13] = 40'b0000000000000000000011111111111111110000;
assign Roles_Image_2[14] = 40'b0000000000000000000011111111111111110000;
assign Roles_Image_2[15] = 40'b1100000000000000001111111111000000000000;
assign Roles_Image_2[16] = 40'b1100000000000000001111111111000000000000;
assign Roles_Image_2[17] = 40'b1100000000000001111111111111000000000000;
assign Roles_Image_2[18] = 40'b1100000000000001111111111111000000000000;
assign Roles_Image_2[19] = 40'b1111000000001111111111111111111100000000;
assign Roles_Image_2[20] = 40'b1111000000001111111111111111111100000000;
assign Roles_Image_2[21] = 40'b1111110000111111111111111111001100000000;
assign Roles_Image_2[22] = 40'b1111110000111111111111111111001100000000;
assign Roles_Image_2[23] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_2[24] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_2[25] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_2[26] = 40'b1111111111111111111111111111000000000000;
assign Roles_Image_2[27] = 40'b0011111111111111111111111111000000000000;
assign Roles_Image_2[28] = 40'b0011111111111111111111111100000000000000;
assign Roles_Image_2[29] = 40'b0000111111111111111111111100000000000000;
assign Roles_Image_2[30] = 40'b0000111111111111111111111100000000000000;
assign Roles_Image_2[31] = 40'b0000001111111111111111110000000000000000;
assign Roles_Image_2[32] = 40'b0000001111111111111111110000000000000000;
assign Roles_Image_2[33] = 40'b0000000011111111111111000000000000000000;
assign Roles_Image_2[34] = 40'b0000000011111111111111000000000000000000;
assign Roles_Image_2[35] = 40'b0000000000111111000011111000000000000000;
assign Roles_Image_2[36] = 40'b0000000000111111000011111000000000000000;
assign Roles_Image_2[37] = 40'b0000000000111100000000000000000000000000;
assign Roles_Image_2[38] = 40'b0000000000111100000000000000000000000000;
assign Roles_Image_2[39] = 40'b0000000000110000000000000000000000000000;
assign Roles_Image_2[40] = 40'b0000000000110000000000000000000000000000;
assign Roles_Image_2[41] = 40'b0000000000111100000000000000000000000000;
assign Roles_Image_2[42] = 40'b0000000000111100000000000000000000000000;


wire [ 0 : 14] Cactus_Image[ 0 : 32];
assign Cactus_Image[0] = 15'b000000111000000;
assign Cactus_Image[1] = 15'b000001111100000;
assign Cactus_Image[2] = 15'b000001111100000;
assign Cactus_Image[3] = 15'b000001111100000;
assign Cactus_Image[4] = 15'b000001111100010;
assign Cactus_Image[5] = 15'b000001111100111;
assign Cactus_Image[6] = 15'b000001111100111;
assign Cactus_Image[7] = 15'b000001111100111;
assign Cactus_Image[8] = 15'b010001111100111;
assign Cactus_Image[9] = 15'b111001111100111;
assign Cactus_Image[10] = 15'b111001111100111;
assign Cactus_Image[11] = 15'b111001111100111;
assign Cactus_Image[12] = 15'b111001111100111;
assign Cactus_Image[13] = 15'b111001111100111;
assign Cactus_Image[14] = 15'b111001111100111;
assign Cactus_Image[15] = 15'b111001111111111;
assign Cactus_Image[16] = 15'b111001111111110;
assign Cactus_Image[17] = 15'b111001111111100;
assign Cactus_Image[18] = 15'b111001111100000;
assign Cactus_Image[19] = 15'b111111111100000;
assign Cactus_Image[20] = 15'b011111111100000;
assign Cactus_Image[21] = 15'b001111111100000;
assign Cactus_Image[22] = 15'b000001111100000;
assign Cactus_Image[23] = 15'b000001111100000;
assign Cactus_Image[24] = 15'b000001111100000;
assign Cactus_Image[25] = 15'b000001111100000;
assign Cactus_Image[26] = 15'b000001111100000;
assign Cactus_Image[27] = 15'b000001111100000;
assign Cactus_Image[28] = 15'b000001111100000;
assign Cactus_Image[29] = 15'b000001111100000;
assign Cactus_Image[30] = 15'b000001111100000;
assign Cactus_Image[31] = 15'b000001111100000;
assign Cactus_Image[32] = 15'b000001111100000;


wire [ 0 : 17] Fire_Image[ 0 : 9];
assign Fire_Image[0] = 18'b110000000000000000;
assign Fire_Image[1] = 18'b111000000111100000;
assign Fire_Image[2] = 18'b111111011111000000;
assign Fire_Image[3] = 18'b111111111111111000;
assign Fire_Image[4] = 18'b111111111111111110;
assign Fire_Image[5] = 18'b011111111111111111;
assign Fire_Image[6] = 18'b011111111111111000;
assign Fire_Image[7] = 18'b001111111111110000;
assign Fire_Image[8] = 18'b000011111111100000;
assign Fire_Image[9] = 18'b000000111111000000;


wire [ 0 : 275] Ranther_Image[ 0 : 85];
assign Ranther_Image[0] = 276'b000000000000000000000000000000001111000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[1] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[2] = 276'b000000000000000000000000011000000000000001100000000000000000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[3] = 276'b000000000000000000000000011000000000000001100000000000000000000001100000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[4] = 276'b000000000000000000000000001000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[5] = 276'b000000000000000000000000010000000000000000000011111111111111110000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[6] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[7] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[8] = 276'b000000000000000000010000110000001100000000000000010000000100000000000000000100000001000010000000000000000000000000000000000000000000000000000000000000000000000001000000010000000100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[9] = 276'b000000000000000000100000011000000110000000000000010000000100000000000000000100000001000001000000000000000000000000000000000000000000000000000000000000000000000001000000010000000100000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[10] = 276'b000000000000000001000000000100000001000000000000010000000100000000000000000100000001000000100000000000000000000000000000000000000000000000000000000000000000000001000000010000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[11] = 276'b000000000000000001000000000000000000000000000000010000000100000000000000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000001000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[12] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000001000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[13] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000001000000010000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[14] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000010000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[15] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000010000000100000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[16] = 276'b000000000000000010000000000000000000000011110000000000000000000011110000010000000100000000010000000000000000000000000000000000000000000000000000111100001111000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[17] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000100000001000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[18] = 276'b000000000000000010000000000000000000000000000000000000000000000000000000100000001000000000010000011000000000000000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[19] = 276'b000000000000000001000000000000000000000000000000000000000000000000000000100000001000000000100000011000000000000000000000000000000110000001100000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[20] = 276'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[21] = 276'b000000000000000000100000000000000000000000000000000000000000000000000000000000000000000001000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[22] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[23] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[24] = 276'b000000000000000000000000110000000011100000000000000000000011100000000000000000001000000000000000000000000000000011000000000000000000000000000000000000000001000000000000000000000000000000000000000000001000000000000000110000000000000000000000000000000000000000000000110000001000;
assign Ranther_Image[25] = 276'b000000000000000000000000011000000100000000000000000000000100000000000000000000000100000000000000000000000000000001100000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000011000000000000000000000000000000000000000000000011000000100;
assign Ranther_Image[26] = 276'b000000000000000000000000000100001000000000000000000000001000000000000000000000000010000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000100000000000000000000000000000000000000000000000100000010;
assign Ranther_Image[27] = 276'b000000000000000000000000000000010000000000000000000000010000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010;
assign Ranther_Image[28] = 276'b000000000000000000000000000000010110000000000000000000010110000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001;
assign Ranther_Image[29] = 276'b000000000000000000000000000000011001000000000000000000011001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001;
assign Ranther_Image[30] = 276'b000000000000000000000000000000010000100000000000000000010000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001;
assign Ranther_Image[31] = 276'b000000000000000000000000000000010000100000000000000000010000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001;
assign Ranther_Image[32] = 276'b000000000000000000000000000000010000100000000000000000010000100000000000000000000001000000000000000000000000000000000000111100000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000001111000000000000000000000000000000000000000000000001;
assign Ranther_Image[33] = 276'b000000000000000000000000000000010000100000000000000000010000100000000000000000000001000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000001;
assign Ranther_Image[34] = 276'b000000000000000000000000000000001001000000000000000000001001000000000000000000000001000000000000000000000000000000000000000000000110000000000000000000001000000000000000000000000000000000000000000000000001000001100000000000000000000001100000000000000000000001100000000000000001;
assign Ranther_Image[35] = 276'b000000000000000000000000000000000110000000000000000000000110000000000000000000000010000000000000000000000000000000000000000000000110000000000000000000000100000000000000000000000000000000000000000000000010000001100000000000000000000001100000000000000000000001100000000000000010;
assign Ranther_Image[36] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010;
assign Ranther_Image[37] = 276'b000000000000000000000000000000000000001111111100000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000100000000000000000000000000000000000011111111111111110000000000000000000100;
assign Ranther_Image[38] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[39] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[40] = 276'b000000000000000000000000000100000000001110111000000000000000000010000000010000000000000000000000000000000000000000000000000000000000000010000000000000000000000011000000000000000000000000000000110000000000000000000000110000001100000000000000000000000000000000000000010000000000;
assign Ranther_Image[41] = 276'b000000000000000000000000001000000000000100010000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000001000000000000000000000001100000000000000000000000000000011000000000000000000000011000000110000000000000000000000000000000000000010000000000;
assign Ranther_Image[42] = 276'b000000000000000000000000010000000000000100010000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000010000000000000000000000000000000100000000000000000000000100000001000000000000000000000000000000000000010000000000;
assign Ranther_Image[43] = 276'b000000000000000000000000010000000000000010100000000000000000000000100000010000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
assign Ranther_Image[44] = 276'b000000000000000000000000100000000000000010100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[45] = 276'b000000000000000000000000100000000000000010100000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[46] = 276'b000000000000000000000000100000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[47] = 276'b000000000000000000000000100000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[48] = 276'b000000000000000000000000100000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000011110000000000000000;
assign Ranther_Image[49] = 276'b000000000000000000000000100000000000000001000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[50] = 276'b000000000000000000000000100000000000000001000000000000000110000000010000000000000000000000000000011000000000000000000000000000000000000000010000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000000000000011000000110000000000000000000000000;
assign Ranther_Image[51] = 276'b000000000000000000000000010000000000000011100000000000000110000000100000000000000000000000000000011000000000000000000000000000000000000000100000000000000000000000000000011000000000000000000000000000000110000000000000000000000000000000000000011000000110000000000000000000000000;
assign Ranther_Image[52] = 276'b000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[53] = 276'b000000000000000000000000001000111111110000000011111111000000000001000000000000000000000000000000000000111111110000000000000000000000000001000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[54] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[55] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[56] = 276'b000000000000000000000000000000001100000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[57] = 276'b000000000000000000000000000000000110000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[58] = 276'b000000000000000000000000000000000001000000000000000000000100000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[59] = 276'b000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000100000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[60] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[61] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[62] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[63] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[64] = 276'b000000000000000000000000000000000000000011110000111100000000000000000000000000000000000011110000000000000100000000000000000000000100000011110000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[65] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[66] = 276'b000000000000000001100000011000000000000000000000000000000000000000000000011000000110000000000000000000001000000000000000000000001000000000000000000000000000000000000000011000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[67] = 276'b000000000000000001100000011000000000000000000000000000000000000000000000011000000110000000000000000000001000000000000000000000001000000000000000000000000000000000000000011000000000000000000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[68] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[69] = 276'b000000111111110000000000000000000000000000000000000000000000001111111100000000000000000000000011111111000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[70] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[71] = 276'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[72] = 276'b000100000010000001100000100000000000000000000000010000000100000000000000000000000001000001100000001000001000000000000000010000000000000000000000000100000001000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[73] = 276'b001000000010000000100000010000000000000000000000010000000100000000000000000000000010000000100000001000000100000000000000010000000000000000000000001000000010000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[74] = 276'b010000000000000000100000001000000000000000000000010000000100000000000000000000000100000000100000000000000010000000000000010000000000000000000000010000000100000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[75] = 276'b010000000010000000100000001000000000000000000000010000000100000000000000000000000100000000100000001000000010000000000000010000000000000000000000010000000100000001000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[76] = 276'b100000000110000000100000000100000000000000000000000000000000000000000000000000001000000000100000011000000001000000000000000000000000000000000000100000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[77] = 276'b100000000010000000100000000100000000000000000000000000000000000000000000000000001000000000100000001000000001000000000000000000000000000000000000100000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[78] = 276'b100000000010000000100000000100000000000000000000000000000000000000000000000000001000000000100000001000000001000000000000000000000000000000000000100000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[79] = 276'b100000000010000000100000000100000000000000000000000000000000000000000000000000001000000000100000001000000001000000000000000000000000000000000000100000001000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[80] = 276'b100000000010000000100000000100000000000011110000000000000000000000000000000000001000000000100000001000000001000000000000000000000000000000000000100000001000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[81] = 276'b100000000010000000100000000100000000000000000000000000000000000000000000000000001000000000100000001000000001000000000000000000000000000000000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[82] = 276'b100000000010000000100000000100000110000000000000000000000000000000000000000000001000000000100000001000000001000001100000000000000000000000000000100000001000000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[83] = 276'b010000000111000001110000001000000110000000000000000000000000000000000000000000000100000001110000011100000010000001100000000000000000000000000000010000000100000001000000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[84] = 276'b010000000000000000000000001000000010000000000000000000000000000000000000000000000100000000000000000000000010000000100000000000000000000000000000010000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
assign Ranther_Image[85] = 276'b001000000000000000000000010000000100000000000000000000000000000000000000000000000010000000000000000000000100000001000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;



/*-------------------------------------------------------*/
endmodule