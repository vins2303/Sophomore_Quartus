library verilog;
use verilog.vl_types.all;
entity cyclonev_fractional_pll is
    generic(
        output_clock_frequency: string  := "";
        reference_clock_frequency: string  := "";
        mimic_fbclk_type: string  := "cdb_pll_mimic_fbclk_gclk";
        dsm_accumulator_reset_value: integer := 0;
        forcelock       : string  := "false";
        nreset_invert   : string  := "false";
        pll_atb         : integer := 0;
        pll_bwctrl      : integer := 10000;
        pll_cmp_buf_dly : string  := "0 ps";
        pll_cp_comp     : string  := "true";
        pll_cp_current  : integer := 20;
        pll_ctrl_override_setting: string  := "false";
        pll_dsm_dither  : string  := "disable";
        pll_dsm_out_sel : string  := "disable";
        pll_dsm_reset   : string  := "false";
        pll_ecn_bypass  : string  := "false";
        pll_ecn_test_en : string  := "false";
        pll_enable      : string  := "true";
        pll_fbclk_mux_1 : string  := "glb";
        pll_fbclk_mux_2 : string  := "fb_1";
        pll_fractional_carry_out: integer := 24;
        pll_fractional_division: integer := 1;
        pll_fractional_division_string: string  := "1";
        pll_fractional_value_ready: string  := "true";
        pll_lf_testen   : string  := "false";
        pll_lock_fltr_cfg: integer := 0;
        pll_lock_fltr_test: string  := "false";
        pll_m_cnt_bypass_en: string  := "false";
        pll_m_cnt_coarse_dly: string  := "0 ps";
        pll_m_cnt_fine_dly: string  := "0 ps";
        pll_m_cnt_hi_div: integer := 1;
        pll_m_cnt_in_src: string  := "ph_mux_clk";
        pll_m_cnt_lo_div: integer := 1;
        pll_m_cnt_odd_div_duty_en: string  := "false";
        pll_m_cnt_ph_mux_prst: integer := 0;
        pll_m_cnt_prst  : integer := 1;
        pll_n_cnt_bypass_en: string  := "false";
        pll_n_cnt_coarse_dly: string  := "0 ps";
        pll_n_cnt_fine_dly: string  := "0 ps";
        pll_n_cnt_hi_div: integer := 1;
        pll_n_cnt_lo_div: integer := 1;
        pll_n_cnt_odd_div_duty_en: string  := "false";
        pll_ref_buf_dly : string  := "0 ps";
        pll_reg_boost   : integer := 0;
        pll_regulator_bypass: string  := "false";
        pll_ripplecap_ctrl: integer := 0;
        pll_slf_rst     : string  := "false";
        pll_tclk_mux_en : string  := "false";
        pll_tclk_sel    : string  := "cdb_pll_tclk_sel_m_src";
        pll_test_enable : string  := "false";
        pll_testdn_enable: string  := "false";
        pll_testup_enable: string  := "false";
        pll_unlock_fltr_cfg: integer := 0;
        pll_vco_div     : integer := 2;
        pll_vco_ph0_en  : string  := "false";
        pll_vco_ph1_en  : string  := "false";
        pll_vco_ph2_en  : string  := "false";
        pll_vco_ph3_en  : string  := "false";
        pll_vco_ph4_en  : string  := "false";
        pll_vco_ph5_en  : string  := "false";
        pll_vco_ph6_en  : string  := "false";
        pll_vco_ph7_en  : string  := "false";
        pll_vctrl_test_voltage: integer := 750;
        vccd0g_atb      : string  := "disable";
        vccd0g_output   : integer := 0;
        vccd1g_atb      : string  := "disable";
        vccd1g_output   : integer := 0;
        vccm1g_tap      : integer := 2;
        vccr_pd         : string  := "false";
        vcodiv_override : string  := "false";
        fractional_pll_index: integer := 1
    );
    port(
        coreclkfb       : in     vl_logic_vector(0 downto 0);
        ecnc1test       : in     vl_logic_vector(0 downto 0);
        ecnc2test       : in     vl_logic_vector(0 downto 0);
        fbclkfpll       : in     vl_logic_vector(0 downto 0);
        lvdsfbin        : in     vl_logic_vector(0 downto 0);
        nresync         : in     vl_logic_vector(0 downto 0);
        pfden           : in     vl_logic_vector(0 downto 0);
        refclkin        : in     vl_logic_vector(0 downto 0);
        shift           : in     vl_logic_vector(0 downto 0);
        shiftdonein     : in     vl_logic_vector(0 downto 0);
        shiften         : in     vl_logic_vector(0 downto 0);
        up              : in     vl_logic_vector(0 downto 0);
        vsspl           : in     vl_logic_vector(0 downto 0);
        zdb             : in     vl_logic_vector(0 downto 0);
        cntnen          : out    vl_logic_vector(0 downto 0);
        fbclk           : out    vl_logic_vector(0 downto 0);
        fblvdsout       : out    vl_logic_vector(0 downto 0);
        lock            : out    vl_logic_vector(0 downto 0);
        mhi             : out    vl_logic_vector(7 downto 0);
        mcntout         : out    vl_logic_vector(0 downto 0);
        plniotribuf     : out    vl_logic_vector(0 downto 0);
        shiftdoneout    : out    vl_logic_vector(0 downto 0);
        tclk            : out    vl_logic_vector(0 downto 0);
        vcoph           : out    vl_logic_vector(7 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of output_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of reference_clock_frequency : constant is 1;
    attribute mti_svvh_generic_type of mimic_fbclk_type : constant is 1;
    attribute mti_svvh_generic_type of dsm_accumulator_reset_value : constant is 1;
    attribute mti_svvh_generic_type of forcelock : constant is 1;
    attribute mti_svvh_generic_type of nreset_invert : constant is 1;
    attribute mti_svvh_generic_type of pll_atb : constant is 1;
    attribute mti_svvh_generic_type of pll_bwctrl : constant is 1;
    attribute mti_svvh_generic_type of pll_cmp_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_comp : constant is 1;
    attribute mti_svvh_generic_type of pll_cp_current : constant is 1;
    attribute mti_svvh_generic_type of pll_ctrl_override_setting : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_dither : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_out_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_dsm_reset : constant is 1;
    attribute mti_svvh_generic_type of pll_ecn_bypass : constant is 1;
    attribute mti_svvh_generic_type of pll_ecn_test_en : constant is 1;
    attribute mti_svvh_generic_type of pll_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_1 : constant is 1;
    attribute mti_svvh_generic_type of pll_fbclk_mux_2 : constant is 1;
    attribute mti_svvh_generic_type of pll_fractional_carry_out : constant is 1;
    attribute mti_svvh_generic_type of pll_fractional_division : constant is 1;
    attribute mti_svvh_generic_type of pll_fractional_division_string : constant is 1;
    attribute mti_svvh_generic_type of pll_fractional_value_ready : constant is 1;
    attribute mti_svvh_generic_type of pll_lf_testen : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_lock_fltr_test : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_hi_div : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_in_src : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_lo_div : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_odd_div_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_ph_mux_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_m_cnt_prst : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_bypass_en : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_coarse_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_fine_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_hi_div : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_lo_div : constant is 1;
    attribute mti_svvh_generic_type of pll_n_cnt_odd_div_duty_en : constant is 1;
    attribute mti_svvh_generic_type of pll_ref_buf_dly : constant is 1;
    attribute mti_svvh_generic_type of pll_reg_boost : constant is 1;
    attribute mti_svvh_generic_type of pll_regulator_bypass : constant is 1;
    attribute mti_svvh_generic_type of pll_ripplecap_ctrl : constant is 1;
    attribute mti_svvh_generic_type of pll_slf_rst : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_mux_en : constant is 1;
    attribute mti_svvh_generic_type of pll_tclk_sel : constant is 1;
    attribute mti_svvh_generic_type of pll_test_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_testdn_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_testup_enable : constant is 1;
    attribute mti_svvh_generic_type of pll_unlock_fltr_cfg : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_div : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph0_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph1_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph2_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph3_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph4_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph5_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph6_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vco_ph7_en : constant is 1;
    attribute mti_svvh_generic_type of pll_vctrl_test_voltage : constant is 1;
    attribute mti_svvh_generic_type of vccd0g_atb : constant is 1;
    attribute mti_svvh_generic_type of vccd0g_output : constant is 1;
    attribute mti_svvh_generic_type of vccd1g_atb : constant is 1;
    attribute mti_svvh_generic_type of vccd1g_output : constant is 1;
    attribute mti_svvh_generic_type of vccm1g_tap : constant is 1;
    attribute mti_svvh_generic_type of vccr_pd : constant is 1;
    attribute mti_svvh_generic_type of vcodiv_override : constant is 1;
    attribute mti_svvh_generic_type of fractional_pll_index : constant is 1;
end cyclonev_fractional_pll;
