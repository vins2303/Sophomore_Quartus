library verilog;
use verilog.vl_types.all;
entity cyclonev_hps_interface_fpga2sdram is
    port(
        cfg_axi_mm_select: in     vl_logic_vector(5 downto 0);
        cfg_cport_rfifo_map: in     vl_logic_vector(17 downto 0);
        cfg_cport_type  : in     vl_logic_vector(11 downto 0);
        cfg_cport_wfifo_map: in     vl_logic_vector(17 downto 0);
        cfg_port_width  : in     vl_logic_vector(11 downto 0);
        cfg_rfifo_cport_map: in     vl_logic_vector(15 downto 0);
        cfg_wfifo_cport_map: in     vl_logic_vector(15 downto 0);
        cmd_data_0      : in     vl_logic_vector(59 downto 0);
        cmd_data_1      : in     vl_logic_vector(59 downto 0);
        cmd_data_2      : in     vl_logic_vector(59 downto 0);
        cmd_data_3      : in     vl_logic_vector(59 downto 0);
        cmd_data_4      : in     vl_logic_vector(59 downto 0);
        cmd_data_5      : in     vl_logic_vector(59 downto 0);
        cmd_port_clk_0  : in     vl_logic;
        cmd_port_clk_1  : in     vl_logic;
        cmd_port_clk_2  : in     vl_logic;
        cmd_port_clk_3  : in     vl_logic;
        cmd_port_clk_4  : in     vl_logic;
        cmd_port_clk_5  : in     vl_logic;
        cmd_valid_0     : in     vl_logic;
        cmd_valid_1     : in     vl_logic;
        cmd_valid_2     : in     vl_logic;
        cmd_valid_3     : in     vl_logic;
        cmd_valid_4     : in     vl_logic;
        cmd_valid_5     : in     vl_logic;
        rd_clk_0        : in     vl_logic;
        rd_clk_1        : in     vl_logic;
        rd_clk_2        : in     vl_logic;
        rd_clk_3        : in     vl_logic;
        rd_ready_0      : in     vl_logic;
        rd_ready_1      : in     vl_logic;
        rd_ready_2      : in     vl_logic;
        rd_ready_3      : in     vl_logic;
        wr_clk_0        : in     vl_logic;
        wr_clk_1        : in     vl_logic;
        wr_clk_2        : in     vl_logic;
        wr_clk_3        : in     vl_logic;
        wr_data_0       : in     vl_logic_vector(89 downto 0);
        wr_data_1       : in     vl_logic_vector(89 downto 0);
        wr_data_2       : in     vl_logic_vector(89 downto 0);
        wr_data_3       : in     vl_logic_vector(89 downto 0);
        wr_valid_0      : in     vl_logic;
        wr_valid_1      : in     vl_logic;
        wr_valid_2      : in     vl_logic;
        wr_valid_3      : in     vl_logic;
        wrack_ready_0   : in     vl_logic;
        wrack_ready_1   : in     vl_logic;
        wrack_ready_2   : in     vl_logic;
        wrack_ready_3   : in     vl_logic;
        wrack_ready_4   : in     vl_logic;
        wrack_ready_5   : in     vl_logic;
        bonding_out_1   : out    vl_logic_vector(3 downto 0);
        bonding_out_2   : out    vl_logic_vector(3 downto 0);
        cmd_ready_0     : out    vl_logic;
        cmd_ready_1     : out    vl_logic;
        cmd_ready_2     : out    vl_logic;
        cmd_ready_3     : out    vl_logic;
        cmd_ready_4     : out    vl_logic;
        cmd_ready_5     : out    vl_logic;
        rd_data_0       : out    vl_logic_vector(79 downto 0);
        rd_data_1       : out    vl_logic_vector(79 downto 0);
        rd_data_2       : out    vl_logic_vector(79 downto 0);
        rd_data_3       : out    vl_logic_vector(79 downto 0);
        rd_valid_0      : out    vl_logic;
        rd_valid_1      : out    vl_logic;
        rd_valid_2      : out    vl_logic;
        rd_valid_3      : out    vl_logic;
        wr_ready_0      : out    vl_logic;
        wr_ready_1      : out    vl_logic;
        wr_ready_2      : out    vl_logic;
        wr_ready_3      : out    vl_logic;
        wrack_data_0    : out    vl_logic_vector(9 downto 0);
        wrack_data_1    : out    vl_logic_vector(9 downto 0);
        wrack_data_2    : out    vl_logic_vector(9 downto 0);
        wrack_data_3    : out    vl_logic_vector(9 downto 0);
        wrack_data_4    : out    vl_logic_vector(9 downto 0);
        wrack_data_5    : out    vl_logic_vector(9 downto 0);
        wrack_valid_0   : out    vl_logic;
        wrack_valid_1   : out    vl_logic;
        wrack_valid_2   : out    vl_logic;
        wrack_valid_3   : out    vl_logic;
        wrack_valid_4   : out    vl_logic;
        wrack_valid_5   : out    vl_logic
    );
end cyclonev_hps_interface_fpga2sdram;
